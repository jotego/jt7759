/*  This file is part of JT7759.
    JT7759 program is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public Licen4se as published by
    the Free Software Foundation, either version 3 of the Licen4se, or
    (at your option) any later version.

    JT7759 program is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public Licen4se for more details.

    You should have received a copy of the GNU General Public Licen4se
    along with JT7759.  If not, see <http://www.gnu.org/licen4ses/>.

    Author: Jose Tejada Gomez. Twitter: @topapate
    Version: 1.0
    Date: 5-7-2020 */

module jt7759_adpcm #(parameter SW=9) (
    input                      rst,
    input                      clk,
    input                      cendec,
    input             [   3:0] encoded,
    output reg signed [SW-1:0] sound
);

// The look-up table could have been compressed. One obvious way is to realize that one
// half of it is just the negative version of the other.
// However, because it will be synthesized as a 1 kilo word memory of 9-bit words, i.e. 1BRAM
// this is the best choice.
// This is generated by the file doc/lut.c

reg  signed [8:0] lut[0:255];
reg  signed [3:0] st_lut[0:7];
reg         [3:0] st;
reg         [3:0] st_delta;
reg  signed [5:0] st_next, st_sum;

function [SW-1:0] sign_ext;
    input signed [8:0] din;
    sign_ext = { {SW-9{din[8]}}, din };
endfunction

always @(*) begin
    st_delta = st_lut[ encoded[2:0] ];
    st_sum   = {2'b0, st } + {{2{st_delta[3]}}, st_delta };
    if( st_sum[5] )
        st_next = 6'd0;
    else if( st_sum[4] )
        st_next = 6'd15;
    else
        st_next = st_sum;
end

always @(posedge clk, posedge rst ) begin
    if( rst ) begin
        sound <= {SW{1'd0}};
        st    <= 4'd0;
    end else if(cendec) begin
        sound <= sound + sign_ext( lut[{st,encoded}] );
        st    <= st_next[3:0];
    end
end

initial begin
    st_lut[0]=-4'd1; st_lut[1]=-4'd1; st_lut[2]=4'd0; st_lut[3]=4'd0;
    st_lut[4]=4'd1;  st_lut[5]=4'd2;  st_lut[6]=4'd2; st_lut[7]=4'd3;
end


initial begin
    lut[8'h00]=9'd0000; lut[8'h01]=9'd0000; lut[8'h02]=9'd0001; lut[8'h03]=9'd0002; 
    lut[8'h04]=9'd0003; lut[8'h05]=9'd0005; lut[8'h06]=9'd0007; lut[8'h07]=9'd0010; 
    lut[8'h08]=9'd0000; lut[8'h09]=9'd0000; lut[8'h0A]=-9'd001; lut[8'h0B]=-9'd002; 
    lut[8'h0C]=-9'd003; lut[8'h0D]=-9'd005; lut[8'h0E]=-9'd007; lut[8'h0F]=-9'd010; 
    lut[8'h10]=9'd0000; lut[8'h11]=9'd0001; lut[8'h12]=9'd0002; lut[8'h13]=9'd0003; 
    lut[8'h14]=9'd0004; lut[8'h15]=9'd0006; lut[8'h16]=9'd0008; lut[8'h17]=9'd0013; 
    lut[8'h18]=9'd0000; lut[8'h19]=-9'd001; lut[8'h1A]=-9'd002; lut[8'h1B]=-9'd003; 
    lut[8'h1C]=-9'd004; lut[8'h1D]=-9'd006; lut[8'h1E]=-9'd008; lut[8'h1F]=-9'd013; 
    lut[8'h20]=9'd0000; lut[8'h21]=9'd0001; lut[8'h22]=9'd0002; lut[8'h23]=9'd0004; 
    lut[8'h24]=9'd0005; lut[8'h25]=9'd0007; lut[8'h26]=9'd0010; lut[8'h27]=9'd0015; 
    lut[8'h28]=9'd0000; lut[8'h29]=-9'd001; lut[8'h2A]=-9'd002; lut[8'h2B]=-9'd004; 
    lut[8'h2C]=-9'd005; lut[8'h2D]=-9'd007; lut[8'h2E]=-9'd010; lut[8'h2F]=-9'd015; 
    lut[8'h30]=9'd0000; lut[8'h31]=9'd0001; lut[8'h32]=9'd0003; lut[8'h33]=9'd0004; 
    lut[8'h34]=9'd0006; lut[8'h35]=9'd0009; lut[8'h36]=9'd0013; lut[8'h37]=9'd0019; 
    lut[8'h38]=9'd0000; lut[8'h39]=-9'd001; lut[8'h3A]=-9'd003; lut[8'h3B]=-9'd004; 
    lut[8'h3C]=-9'd006; lut[8'h3D]=-9'd009; lut[8'h3E]=-9'd013; lut[8'h3F]=-9'd019; 
    lut[8'h40]=9'd0000; lut[8'h41]=9'd0002; lut[8'h42]=9'd0003; lut[8'h43]=9'd0005; 
    lut[8'h44]=9'd0008; lut[8'h45]=9'd0011; lut[8'h46]=9'd0015; lut[8'h47]=9'd0023; 
    lut[8'h48]=9'd0000; lut[8'h49]=-9'd002; lut[8'h4A]=-9'd003; lut[8'h4B]=-9'd005; 
    lut[8'h4C]=-9'd008; lut[8'h4D]=-9'd011; lut[8'h4E]=-9'd015; lut[8'h4F]=-9'd023; 
    lut[8'h50]=9'd0000; lut[8'h51]=9'd0002; lut[8'h52]=9'd0004; lut[8'h53]=9'd0007; 
    lut[8'h54]=9'd0010; lut[8'h55]=9'd0014; lut[8'h56]=9'd0019; lut[8'h57]=9'd0029; 
    lut[8'h58]=9'd0000; lut[8'h59]=-9'd002; lut[8'h5A]=-9'd004; lut[8'h5B]=-9'd007; 
    lut[8'h5C]=-9'd010; lut[8'h5D]=-9'd014; lut[8'h5E]=-9'd019; lut[8'h5F]=-9'd029; 
    lut[8'h60]=9'd0000; lut[8'h61]=9'd0003; lut[8'h62]=9'd0005; lut[8'h63]=9'd0008; 
    lut[8'h64]=9'd0012; lut[8'h65]=9'd0016; lut[8'h66]=9'd0022; lut[8'h67]=9'd0033; 
    lut[8'h68]=9'd0000; lut[8'h69]=-9'd003; lut[8'h6A]=-9'd005; lut[8'h6B]=-9'd008; 
    lut[8'h6C]=-9'd012; lut[8'h6D]=-9'd016; lut[8'h6E]=-9'd022; lut[8'h6F]=-9'd033; 
    lut[8'h70]=9'd0001; lut[8'h71]=9'd0004; lut[8'h72]=9'd0007; lut[8'h73]=9'd0010; 
    lut[8'h74]=9'd0015; lut[8'h75]=9'd0020; lut[8'h76]=9'd0029; lut[8'h77]=9'd0043; 
    lut[8'h78]=-9'd001; lut[8'h79]=-9'd004; lut[8'h7A]=-9'd007; lut[8'h7B]=-9'd010; 
    lut[8'h7C]=-9'd015; lut[8'h7D]=-9'd020; lut[8'h7E]=-9'd029; lut[8'h7F]=-9'd043; 
    lut[8'h80]=9'd0001; lut[8'h81]=9'd0004; lut[8'h82]=9'd0008; lut[8'h83]=9'd0013; 
    lut[8'h84]=9'd0018; lut[8'h85]=9'd0025; lut[8'h86]=9'd0035; lut[8'h87]=9'd0053; 
    lut[8'h88]=-9'd001; lut[8'h89]=-9'd004; lut[8'h8A]=-9'd008; lut[8'h8B]=-9'd013; 
    lut[8'h8C]=-9'd018; lut[8'h8D]=-9'd025; lut[8'h8E]=-9'd035; lut[8'h8F]=-9'd053; 
    lut[8'h90]=9'd0001; lut[8'h91]=9'd0006; lut[8'h92]=9'd0010; lut[8'h93]=9'd0016; 
    lut[8'h94]=9'd0022; lut[8'h95]=9'd0031; lut[8'h96]=9'd0043; lut[8'h97]=9'd0064; 
    lut[8'h98]=-9'd001; lut[8'h99]=-9'd006; lut[8'h9A]=-9'd010; lut[8'h9B]=-9'd016; 
    lut[8'h9C]=-9'd022; lut[8'h9D]=-9'd031; lut[8'h9E]=-9'd043; lut[8'h9F]=-9'd064; 
    lut[8'hA0]=9'd0002; lut[8'hA1]=9'd0007; lut[8'hA2]=9'd0012; lut[8'hA3]=9'd0019; 
    lut[8'hA4]=9'd0027; lut[8'hA5]=9'd0037; lut[8'hA6]=9'd0051; lut[8'hA7]=9'd0076; 
    lut[8'hA8]=-9'd002; lut[8'hA9]=-9'd007; lut[8'hAA]=-9'd012; lut[8'hAB]=-9'd019; 
    lut[8'hAC]=-9'd027; lut[8'hAD]=-9'd037; lut[8'hAE]=-9'd051; lut[8'hAF]=-9'd076; 
    lut[8'hB0]=9'd0002; lut[8'hB1]=9'd0009; lut[8'hB2]=9'd0016; lut[8'hB3]=9'd0024; 
    lut[8'hB4]=9'd0034; lut[8'hB5]=9'd0046; lut[8'hB6]=9'd0064; lut[8'hB7]=9'd0096; 
    lut[8'hB8]=-9'd002; lut[8'hB9]=-9'd009; lut[8'hBA]=-9'd016; lut[8'hBB]=-9'd024; 
    lut[8'hBC]=-9'd034; lut[8'hBD]=-9'd046; lut[8'hBE]=-9'd064; lut[8'hBF]=-9'd096; 
    lut[8'hC0]=9'd0003; lut[8'hC1]=9'd0011; lut[8'hC2]=9'd0019; lut[8'hC3]=9'd0029; 
    lut[8'hC4]=9'd0041; lut[8'hC5]=9'd0057; lut[8'hC6]=9'd0079; lut[8'hC7]=9'd0117; 
    lut[8'hC8]=-9'd003; lut[8'hC9]=-9'd011; lut[8'hCA]=-9'd019; lut[8'hCB]=-9'd029; 
    lut[8'hCC]=-9'd041; lut[8'hCD]=-9'd057; lut[8'hCE]=-9'd079; lut[8'hCF]=-9'd117; 
    lut[8'hD0]=9'd0004; lut[8'hD1]=9'd0013; lut[8'hD2]=9'd0024; lut[8'hD3]=9'd0036; 
    lut[8'hD4]=9'd0050; lut[8'hD5]=9'd0069; lut[8'hD6]=9'd0096; lut[8'hD7]=9'd0143; 
    lut[8'hD8]=-9'd004; lut[8'hD9]=-9'd013; lut[8'hDA]=-9'd024; lut[8'hDB]=-9'd036; 
    lut[8'hDC]=-9'd050; lut[8'hDD]=-9'd069; lut[8'hDE]=-9'd096; lut[8'hDF]=-9'd143; 
    lut[8'hE0]=9'd0004; lut[8'hE1]=9'd0016; lut[8'hE2]=9'd0029; lut[8'hE3]=9'd0044; 
    lut[8'hE4]=9'd0062; lut[8'hE5]=9'd0085; lut[8'hE6]=9'd0118; lut[8'hE7]=9'd0175; 
    lut[8'hE8]=-9'd004; lut[8'hE9]=-9'd016; lut[8'hEA]=-9'd029; lut[8'hEB]=-9'd044; 
    lut[8'hEC]=-9'd062; lut[8'hED]=-9'd085; lut[8'hEE]=-9'd118; lut[8'hEF]=-9'd175; 
    lut[8'hF0]=9'd0006; lut[8'hF1]=9'd0020; lut[8'hF2]=9'd0036; lut[8'hF3]=9'd0054; 
    lut[8'hF4]=9'd0076; lut[8'hF5]=9'd0104; lut[8'hF6]=9'd0144; lut[8'hF7]=9'd0214; 
    lut[8'hF8]=-9'd006; lut[8'hF9]=-9'd020; lut[8'hFA]=-9'd036; lut[8'hFB]=-9'd054; 
    lut[8'hFC]=-9'd076; lut[8'hFD]=-9'd104; lut[8'hFE]=-9'd144; lut[8'hFF]=-9'd214; 
end

endmodule