/*  This file is part of JT7759.
    JT7759 program is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public Licen4se as published by
    the Free Software Foundation, either version 3 of the Licen4se, or
    (at your option) any later version.

    JT7759 program is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public Licen4se for more details.

    You should have received a copy of the GNU General Public Licen4se
    along with JT7759.  If not, see <http://www.gnu.org/licen4ses/>.

    Author: Jose Tejada Gomez. Twitter: @topapate
    Version: 1.0
    Date: 5-7-2020 */

module jt7759_adpcm #(parameter SW=9) (
    input                      rst,
    input                      clk,
    input                      cen_dec,
    input             [   3:0] encoded,
    output reg signed [SW-1:0] sound
);

// The look-up table could have been compressed. One obvious way is to realize that one
// half of it is just the negative version of the other.
// However, because it will be synthesized as a 1 kilo word memory of 9-bit words, i.e. 1BRAM
// this is the best choice.
// This is generated by the file doc/lut.c

reg  signed [8:0] lut[0:255];
reg  signed [3:0] st_lut[0:7];
reg         [3:0] st;
reg         [3:0] st_delta;
reg  signed [5:0] st_next, st_sum;
reg  signed [SW:0] next_snd, lut_step;

function [SW:0] sign_ext;
    input signed [8:0] din;
    sign_ext = { {SW-8{din[8]}}, din };
endfunction

always @(*) begin
    st_delta = st_lut[ encoded[2:0] ];
    st_sum   = {2'b0, st } + {{2{st_delta[3]}}, st_delta };
    if( st_sum[5] )
        st_next = 6'd0;
    else if( st_sum[4] )
        st_next = 6'd15;
    else
        st_next = st_sum;
    lut_step = sign_ext( lut[{st,encoded}] );
    next_snd = { sound[SW-1], sound } + lut_step;
end

always @(posedge clk, posedge rst ) begin
    if( rst ) begin
        sound <= {SW{1'd0}};
        st    <= 4'd0;
    end else if(cen_dec) begin
        if( next_snd[SW]==next_snd[SW-1] )
            sound <= next_snd[SW-1:0];
        else sound <= next_snd[SW] ? {1'b1,{SW-1{1'b0}}} : {1'b0,{SW-1{1'b1}}};
        st    <= st_next[3:0];
    end
end

initial begin
    st_lut[0]=-4'd1; st_lut[1]=-4'd1; st_lut[2]=4'd0; st_lut[3]=4'd0;
    st_lut[4]=4'd1;  st_lut[5]=4'd2;  st_lut[6]=4'd2; st_lut[7]=4'd3;
end


initial begin
    lut[8'h00]= 8'd0;  lut[8'h01]= 8'd0;   lut[8'h02]= 8'd1;   lut[8'h03]= 8'd2;
    lut[8'h04]= 8'd3;  lut[8'h05]= 8'd5;   lut[8'h06]= 8'd7;   lut[8'h07]= 8'd10;
    lut[8'h08]= 8'd0;  lut[8'h09]= 8'd0;   lut[8'h0A]=-8'd1;   lut[8'h0B]=-8'd2;
    lut[8'h0C]=-8'd3;  lut[8'h0D]=-8'd5;   lut[8'h0E]=-8'd7;   lut[8'h0F]=-8'd10;
    lut[8'h10]= 8'd0;  lut[8'h11]= 8'd1;   lut[8'h12]= 8'd2;   lut[8'h13]= 8'd3;
    lut[8'h14]= 8'd4;  lut[8'h15]= 8'd6;   lut[8'h16]= 8'd8;   lut[8'h17]= 8'd13;
    lut[8'h18]= 8'd0;  lut[8'h19]=-8'd1;   lut[8'h1A]=-8'd2;   lut[8'h1B]=-8'd3;
    lut[8'h1C]=-8'd4;  lut[8'h1D]=-8'd6;   lut[8'h1E]=-8'd8;   lut[8'h1F]=-8'd13;
    lut[8'h20]= 8'd0;  lut[8'h21]= 8'd1;   lut[8'h22]= 8'd2;   lut[8'h23]= 8'd4;
    lut[8'h24]= 8'd5;  lut[8'h25]= 8'd7;   lut[8'h26]= 8'd10;  lut[8'h27]= 8'd15;
    lut[8'h28]= 8'd0;  lut[8'h29]=-8'd1;   lut[8'h2A]=-8'd2;   lut[8'h2B]=-8'd4;
    lut[8'h2C]=-8'd5;  lut[8'h2D]=-8'd7;   lut[8'h2E]=-8'd10;  lut[8'h2F]=-8'd15;
    lut[8'h30]= 8'd0;  lut[8'h31]= 8'd1;   lut[8'h32]= 8'd3;   lut[8'h33]= 8'd4;
    lut[8'h34]= 8'd6;  lut[8'h35]= 8'd9;   lut[8'h36]= 8'd13;  lut[8'h37]= 8'd19;
    lut[8'h38]= 8'd0;  lut[8'h39]=-8'd1;   lut[8'h3A]=-8'd3;   lut[8'h3B]=-8'd4;
    lut[8'h3C]=-8'd6;  lut[8'h3D]=-8'd9;   lut[8'h3E]=-8'd13;  lut[8'h3F]=-8'd19;
    lut[8'h40]= 8'd0;  lut[8'h41]= 8'd2;   lut[8'h42]= 8'd3;   lut[8'h43]= 8'd5;
    lut[8'h44]= 8'd8;  lut[8'h45]= 8'd11;  lut[8'h46]= 8'd15;  lut[8'h47]= 8'd23;
    lut[8'h48]= 8'd0;  lut[8'h49]=-8'd2;   lut[8'h4A]=-8'd3;   lut[8'h4B]=-8'd5;
    lut[8'h4C]=-8'd8;  lut[8'h4D]=-8'd11;  lut[8'h4E]=-8'd15;  lut[8'h4F]=-8'd23;
    lut[8'h50]= 8'd0;  lut[8'h51]= 8'd2;   lut[8'h52]= 8'd4;   lut[8'h53]= 8'd7;
    lut[8'h54]= 8'd10; lut[8'h55]= 8'd14;  lut[8'h56]= 8'd19;  lut[8'h57]= 8'd29;
    lut[8'h58]= 8'd0;  lut[8'h59]=-8'd2;   lut[8'h5A]=-8'd4;   lut[8'h5B]=-8'd7;
    lut[8'h5C]=-8'd10; lut[8'h5D]=-8'd14;  lut[8'h5E]=-8'd19;  lut[8'h5F]=-8'd29;
    lut[8'h60]= 8'd0;  lut[8'h61]= 8'd3;   lut[8'h62]= 8'd5;   lut[8'h63]= 8'd8;
    lut[8'h64]= 8'd12; lut[8'h65]= 8'd16;  lut[8'h66]= 8'd22;  lut[8'h67]= 8'd33;
    lut[8'h68]= 8'd0;  lut[8'h69]=-8'd3;   lut[8'h6A]=-8'd5;   lut[8'h6B]=-8'd8;
    lut[8'h6C]=-8'd12; lut[8'h6D]=-8'd16;  lut[8'h6E]=-8'd22;  lut[8'h6F]=-8'd33;
    lut[8'h70]= 8'd1;  lut[8'h71]= 8'd4;   lut[8'h72]= 8'd7;   lut[8'h73]= 8'd10;
    lut[8'h74]= 8'd15; lut[8'h75]= 8'd20;  lut[8'h76]= 8'd29;  lut[8'h77]= 8'd43;
    lut[8'h78]=-8'd1;  lut[8'h79]=-8'd4;   lut[8'h7A]=-8'd7;   lut[8'h7B]=-8'd10;
    lut[8'h7C]=-8'd15; lut[8'h7D]=-8'd20;  lut[8'h7E]=-8'd29;  lut[8'h7F]=-8'd43;
    lut[8'h80]= 8'd1;  lut[8'h81]= 8'd4;   lut[8'h82]= 8'd8;   lut[8'h83]= 8'd13;
    lut[8'h84]= 8'd18; lut[8'h85]= 8'd25;  lut[8'h86]= 8'd35;  lut[8'h87]= 8'd53;
    lut[8'h88]=-8'd1;  lut[8'h89]=-8'd4;   lut[8'h8A]=-8'd8;   lut[8'h8B]=-8'd13;
    lut[8'h8C]=-8'd18; lut[8'h8D]=-8'd25;  lut[8'h8E]=-8'd35;  lut[8'h8F]=-8'd53;
    lut[8'h90]= 8'd1;  lut[8'h91]= 8'd6;   lut[8'h92]= 8'd10;  lut[8'h93]= 8'd16;
    lut[8'h94]= 8'd22; lut[8'h95]= 8'd31;  lut[8'h96]= 8'd43;  lut[8'h97]= 8'd64;
    lut[8'h98]=-8'd1;  lut[8'h99]=-8'd6;   lut[8'h9A]=-8'd10;  lut[8'h9B]=-8'd16;
    lut[8'h9C]=-8'd22; lut[8'h9D]=-8'd31;  lut[8'h9E]=-8'd43;  lut[8'h9F]=-8'd64;
    lut[8'hA0]= 8'd2;  lut[8'hA1]= 8'd7;   lut[8'hA2]= 8'd12;  lut[8'hA3]= 8'd19;
    lut[8'hA4]= 8'd27; lut[8'hA5]= 8'd37;  lut[8'hA6]= 8'd51;  lut[8'hA7]= 8'd76;
    lut[8'hA8]=-8'd2;  lut[8'hA9]=-8'd7;   lut[8'hAA]=-8'd12;  lut[8'hAB]=-8'd19;
    lut[8'hAC]=-8'd27; lut[8'hAD]=-8'd37;  lut[8'hAE]=-8'd51;  lut[8'hAF]=-8'd76;
    lut[8'hB0]= 8'd2;  lut[8'hB1]= 8'd9;   lut[8'hB2]= 8'd16;  lut[8'hB3]= 8'd24;
    lut[8'hB4]= 8'd34; lut[8'hB5]= 8'd46;  lut[8'hB6]= 8'd64;  lut[8'hB7]= 8'd96;
    lut[8'hB8]=-8'd2;  lut[8'hB9]=-8'd9;   lut[8'hBA]=-8'd16;  lut[8'hBB]=-8'd24;
    lut[8'hBC]=-8'd34; lut[8'hBD]=-8'd46;  lut[8'hBE]=-8'd64;  lut[8'hBF]=-8'd96;
    lut[8'hC0]= 8'd3;  lut[8'hC1]= 8'd11;  lut[8'hC2]= 8'd19;  lut[8'hC3]= 8'd29;
    lut[8'hC4]= 8'd41; lut[8'hC5]= 8'd57;  lut[8'hC6]= 8'd79;  lut[8'hC7]= 8'd117;
    lut[8'hC8]=-8'd3;  lut[8'hC9]=-8'd11;  lut[8'hCA]=-8'd19;  lut[8'hCB]=-8'd29;
    lut[8'hCC]=-8'd41; lut[8'hCD]=-8'd57;  lut[8'hCE]=-8'd79;  lut[8'hCF]=-8'd117;
    lut[8'hD0]= 8'd4;  lut[8'hD1]= 8'd13;  lut[8'hD2]= 8'd24;  lut[8'hD3]= 8'd36;
    lut[8'hD4]= 8'd50; lut[8'hD5]= 8'd69;  lut[8'hD6]= 8'd96;  lut[8'hD7]= 8'd143;
    lut[8'hD8]=-8'd4;  lut[8'hD9]=-8'd13;  lut[8'hDA]=-8'd24;  lut[8'hDB]=-8'd36;
    lut[8'hDC]=-8'd50; lut[8'hDD]=-8'd69;  lut[8'hDE]=-8'd96;  lut[8'hDF]=-8'd143;
    lut[8'hE0]= 8'd4;  lut[8'hE1]= 8'd16;  lut[8'hE2]= 8'd29;  lut[8'hE3]= 8'd44;
    lut[8'hE4]= 8'd62; lut[8'hE5]= 8'd85;  lut[8'hE6]= 8'd118; lut[8'hE7]= 8'd175;
    lut[8'hE8]=-8'd4;  lut[8'hE9]=-8'd16;  lut[8'hEA]=-8'd29;  lut[8'hEB]=-8'd44;
    lut[8'hEC]=-8'd62; lut[8'hED]=-8'd85;  lut[8'hEE]=-8'd118; lut[8'hEF]=-8'd175;
    lut[8'hF0]= 8'd6;  lut[8'hF1]= 8'd20;  lut[8'hF2]= 8'd36;  lut[8'hF3]= 8'd54;
    lut[8'hF4]= 8'd76; lut[8'hF5]= 8'd104; lut[8'hF6]= 8'd144; lut[8'hF7]= 8'd214;
    lut[8'hF8]=-8'd6;  lut[8'hF9]=-8'd20;  lut[8'hFA]=-8'd36;  lut[8'hFB]=-8'd54;
    lut[8'hFC]=-8'd76; lut[8'hFD]=-8'd104; lut[8'hFE]=-8'd144; lut[8'hFF]=-8'd214;
end

endmodule